library ieee;

use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library nigella;

package constants is 

	constant prog_mem_addr_top : integer = 65535;
		
end package;
		